module and_gate_st(input A, input B, output Y); 
	assign Y = A&B;
endmodule
